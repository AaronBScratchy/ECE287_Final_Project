module frogger(
	input clock,     
    input reset,     
    output wire hsync,    // HSYNC (to VGA connector)
    output wire vsync,    // VSYNC (to VGA connctor)
    output [7:0] red,     // RED (to resistor DAC VGA connector)
    output [7:0] green,   // GREEN (to resistor DAC to VGA connector)
    output [7:0] blue,    // BLUE (to resistor DAC to VGA connector)
    output sync,          // SYNC to VGA connector
    output clk,           // CLK to VGA connector
    output blank          // BLANK to VGA connector
);

reg [7:0]color_in;

wire clk_25M;
Clock_divider my_25_MHz(clock, clk_25M);

/*
input wire clock,     // 25 MHz
    input wire reset,     // Active high
    input [7:0] color_in, // Pixel color data (RRRGGGBB)
    output [9:0] next_x,  // x-coordinate of NEXT pixel that will be drawn
    output [9:0] next_y,  // y-coordinate of NEXT pixel that will be drawn
    output wire hsync,    // HSYNC (to VGA connector)
    output wire vsync,    // VSYNC (to VGA connctor)
    output [7:0] red,     // RED (to resistor DAC VGA connector)
    output [7:0] green,   // GREEN (to resistor DAC to VGA connector)
    output [7:0] blue,    // BLUE (to resistor DAC to VGA connector)
    output sync,          // SYNC to VGA connector
    output clk,           // CLK to VGA connector
    output blank          // BLANK to VGA connector
*/

wire next_x;
wire next_y;

vga_driver my_vga_driver(clk_25M, reset, color_in, next_x, next_y, hsync, vsync, red, green, blue, sync, clk, blank);

always @(posedge clk_25M) begin
	if(next_y < 10'd20) begin
		color_in <= 8'b11100000;
	end
	else begin
		color_in <= 8'b00000000;
	end
end

endmodule
